// Copyright 2025 Maktab-e-Digital Systems Lahore.
// Licensed under the Apache License, Version 2.0, see LICENSE file for details.
// SPDX-License-Identifier: Apache-2.0
// Description : This file contains the test bench for the modular testing of 4 way set associative cache memory.
// Author:  Eman Nasarrr.
// Date: 10th, August, 2025.
// ADD FILE HERE
