// ADD FILE HERE
